module ();
input ;
output ;

endmodule

/*
module endmodule 
assign wire reg
begin end 
initial always
function endfunction 
task endtask
case default endcase
parameter 
posedge negedge
*/